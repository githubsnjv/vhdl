`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:11:13 02/09/2022 
// Design Name: 
// Module Name:    ripplefulladder_design_sanjeev 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module ripplefulladder_design_sanjeev(
    input p,
    input q,
    input r,
    output sr,
    output cr
    );


endmodule
