`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:17:29 02/09/2022 
// Design Name: 
// Module Name:    fourbitadder_design_sanjeev 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module fourbitadder_design_sanjeev(
    input a,
    input b,
    input c,
    output sum4,
    output carry4
    );


endmodule
