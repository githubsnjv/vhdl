`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:20:44 02/09/2022 
// Design Name: 
// Module Name:    decoder_design_sanjeev 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module decoder_design_sanjeev(
    input a1,
    input a0,
    input e,
    output y3,
    output y2,
    input y1,
    output y0
    );


endmodule
